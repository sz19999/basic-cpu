// ALU module

module alu();



endmodule
// top module

module top(clk, Din, run, resetn, done, bus_out, registers, counter_out);

parameter word = 16;
parameter r = 8;

input [word-1:0] Din;
input clk, run, resetn;
output done;
output [word-1:0] bus_out;
output [word*r-1:0] registers;	// [R7, ..., R0]
output [1:0] counter_out;

wire clear;
wire IRin, Ain, Gin;
wire DINout, Gout;
wire [7:0] Rout, Rin;
wire [word-1:0] IR, bus ,R_0, R_1, R_2, R_3, R_4, R_5, R_6, R_7, G_to_mux, alu_to_G, A_to_alu;
wire [8:0] IR_to_control;
wire [1:0] alu_op;
wire [1:0] counter;

assign registers = {R_7, R_6, R_5, R_4, R_3, R_2, R_1, R_0},
		 bus_out = bus,
		 IR_to_control = IR[8:0],
		 counter_out = counter;
		 
// counter
counter counter1 (
	.clk(clk),
	.clear(clear),
	.count(counter) 
);

// control unit
control_unit control_unit1 (
    .run(run),
	 .resetn(resetn),
	 .IR(IR_to_control),
	 .counter(counter),
	 .clear(clear),
	 .IRin(IRin),
	 .DINout(DINout),
	 .Rout(Rout),
	 .Gout(Gout),
	 .Rin(Rin),
	 .Gin(Gin),
	 .Ain(Ain),
	 .alu_op(alu_op), 
	 .done(done)
);

// mux
mux4x16 mux1 (
	.din(Din),
	.registers({G_to_mux, R_7, R_6, R_5, R_4, R_3, R_2, R_1, R_0}),
	.select({Rout, Gout, DINout}),
	.bus(bus)
);

// ALU
alu alu1 (
	.alu_op(alu_op),
	.A(A_to_alu),
	.bus(bus),
	.G(alu_to_G)
);

// registers
reg16 IR1 (
	.clk(clk),
	.load(IRin),
	.vecin(Din),
	.vecout(IR)
);

reg16 R0 (
	.clk(clk),
	.load(Rin[0]),
	.vecin(bus),
	.vecout(R_0)
);

reg16 R1 (
	.clk(clk),
	.load(Rin[1]),
	.vecin(bus),
	.vecout(R_1)
);

reg16 R2 (
	.clk(clk),
	.load(Rin[2]),
	.vecin(bus),
	.vecout(R_2)
);

reg16 R3 (
	.clk(clk),
	.load(Rin[3]),
	.vecin(bus),
	.vecout(R_3)
);

reg16 R4 (
	.clk(clk),
	.load(Rin[4]),
	.vecin(bus),
	.vecout(R_4)
);

reg16 R5 (
	.clk(clk),
	.load(Rin[5]),
	.vecin(bus),
	.vecout(R_5)
);

reg16 R6 (
	.clk(clk),
	.load(Rin[6]),
	.vecin(bus),
	.vecout(R_6)
);

reg16 R7 (
	.clk(clk),
	.load(Rin[7]),
	.vecin(bus),
	.vecout(R_7)
);


reg16 A (
	.clk(clk),
	.load(Ain),
	.vecin(bus),
	.vecout(A_to_alu)
);

reg16 G (
	.clk(clk),
	.load(Gin),
	.vecin(alu_to_G),
	.vecout(G_to_mux)
);

endmodule
// top module

module top();



endmodule